/*
 * Copyright (c) 2024 Drago Markov
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module tt_um_adder4 (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

  // All output pins must be assigned. If not used, assign to 0.
    assign uo_out[6:4] = 0;  // Example: ou_out is the sum of ui_in and uio_in
    assign uio_out = 0;
  assign uio_oe  = 0;
  adder4 tt_um_adder4(
      .A (ui_in[3:0]),
      .B (ui_in[7:4]),
      .S (uo_out[3:0]),
      .C4 (uo_out[7])
  );
    
endmodule
